// !!! order is important
package spi_dv_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "spi_seq_item.sv"
    `include "spi_seq_lib.sv"
    `include "spi_seqr_base.sv"
    `include "spi_driver.sv"
    `include "spi_monitor.sv"
    `include "spi_agent_base.sv"
    `include "spi_scoreboard.sv"
    `include "spi_master_env_base.sv"
    `include "spi_master_test.sv"

endpackage