class spi_master_test extends uvm_test;
    `uvm_component_utils (spi_master_test);

    
    function new();
        
    endfunction //new()
endclass //spi_master_test